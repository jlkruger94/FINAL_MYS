constant rom : integer_array := (18,
-12,
67,
-46,
90,
-23,
50,
40,
-5,
58,
5,
-2,
34,
-38,
-12,
-8,
-78,
-17,
-50,
-86,
1,
-69,
-38,
49,
-52,
72,
107,
-8,
234,
114,
38,
507,
-291,
741,
-291,
507,
38,
114,
234,
-8,
107,
72,
-52,
49,
-38,
-69,
1,
-86,
-50,
-17,
-78,
-8,
-12,
-38,
34,
-2,
5,
58,
-5,
40,
50,
-23,
90,
-46,
67,
-12,
18
);